`ifndef ASSERT
`define ASSERT

module axi_assertion();
endmodule

`endif
